package i2s_transmitter_pkg;

typedef enum logic [1:0] {IDLE, LOAD, TRANSMIT} state_t;

endpackage