package T_bird_tail_light_FSM_pkg;

    typedef enum bit [2:0] {IDLE, L1, L2, L3, LR3, R1, R2, R3} state_t;
    
endpackage