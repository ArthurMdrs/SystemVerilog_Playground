localparam int WIDTH = 8;
localparam int STAGES = 5;
localparam int RATE = 16;
localparam bit DnI = 0;
