localparam int WIDTH = 8;
localparam int STAGES = 3;
localparam int RATE = 8;
localparam bit DnI = 1;
