localparam int WIDTH = 8;
localparam int STAGES = 6;
localparam int RATE = 8;
